module CommTB ();



endmodule