module saturate_tb ();

endmodule