module UART_wrapper ();

endmodule