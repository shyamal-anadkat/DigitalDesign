module synth_detect(asynth_sig_in, clk, fall_edge);

input asynth_sig_in;
input clk;
output fall_edge;


endmodule
