module ringosc(clk, rst, en, r_out);

input clk, rst;
input en;
output r_out;




endmodule
